module ram8 (out, in, address, clk);
	output [15:0] out;
	input [15:0] in; input [15:0] address; input clk;
