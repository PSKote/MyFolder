module alu (out, zr, ng, c ,x, y);
	output [15:0] out; output zr, ng;
	input [15:0] x ; input [15:0] y ; 
	input [5:0]c ;
	

endmodule 
